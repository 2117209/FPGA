//***************************************************************/
//模块名: mux21
//作 者: Hang Liu

//用 途：多路选择器，用于选择立即数还是数据；
//版本说明:
//***************************************************************/
module mux21 (
    input sel,
    input [7:0] in1,in2,
    output [7:0] out
);
assign out=sel?in2:in1;

endmodule //mux21